module <name>_tb; 
  reg <input>;
  wire <output>

  <module_name> uut();

  initial begin
     $dumpfile("<waveform_file>.vcd");
     $dumpvars();

  end 
endmodule
