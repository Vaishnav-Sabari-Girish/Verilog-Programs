module <name> {

};

endmodule
